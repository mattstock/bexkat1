module mem_select(address, flash, dram, sram0, sram1, led_matrix, monitor, kbd, encoder, serial0, serial1, serial2, switch, spi, invalid);

input [31:0] address;
output flash;
output dram;
output sram0;
output sram1;
output monitor;
output led_matrix;
output kbd;
output encoder;
output serial0;
output serial1;
output serial2;
output invalid;
output switch;
output spi;

// Simple memory map for now
assign monitor =     (address >= 'hffc00000);
assign led_matrix =  (address >= 'hff410000 && address <= 'hff4113ff);
assign spi =         (address >= 'hff400060 && address <= 'hff40006f);
assign serial2 =     (address >= 'hff400050 && address <= 'hff40005f);
assign switch =      (address >= 'hff400040 && address <= 'hff40004f);
assign kbd =         (address >= 'hff400030 && address <= 'hff40003f);
assign serial1 =     (address >= 'hff400020 && address <= 'hff40002f);
assign serial0 =     (address >= 'hff400010 && address <= 'hff40001f);
assign encoder =     (address >= 'hff400000 && address <= 'hff40000f);
assign flash =       (address >= 'hfe000000 && address <= 'hfe3fffff);
assign dram = 1'b0;
assign sram1 =       (address >= 'h00080000 && address <= 'h000fffff);
assign sram0 =       (address >= 'h00000000 && address <= 'h0007ffff);
assign invalid = ~|{monitor, led_matrix, kbd, serial0, serial1, serial2, spi, encoder, flash, dram, sram0, sram1, switch};
endmodule
