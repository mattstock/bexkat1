// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: shift.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 16.1.0 Build 196 10/24/2016 SJ Lite Edition
// ************************************************************


//Copyright (C) 2016  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module shift (
	aclr,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps1x,
	taps2x,
	taps3x,
	taps4x);

	input	  aclr;
	input	  clock;
	input	[160:0]  shiftin;
	output	[160:0]  shiftout;
	output	[160:0]  taps0x;
	output	[160:0]  taps1x;
	output	[160:0]  taps2x;
	output	[160:0]  taps3x;
	output	[160:0]  taps4x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  aclr;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [160:0] sub_wire0;
	wire [804:0] sub_wire1;
	wire [160:0] shiftout = sub_wire0[160:0];
	wire [804:644] sub_wire9 = sub_wire1[804:644];
	wire [643:483] sub_wire8 = sub_wire1[643:483];
	wire [643:483] sub_wire7 = sub_wire8[643:483];
	wire [482:322] sub_wire6 = sub_wire1[482:322];
	wire [482:322] sub_wire5 = sub_wire6[482:322];
	wire [321:161] sub_wire4 = sub_wire1[321:161];
	wire [321:161] sub_wire3 = sub_wire4[321:161];
	wire [160:0] sub_wire2 = sub_wire1[160:0];
	wire [160:0] taps0x = sub_wire2[160:0];
	wire [160:0] taps1x = sub_wire3[321:161];
	wire [160:0] taps2x = sub_wire5[482:322];
	wire [160:0] taps3x = sub_wire7[643:483];
	wire [160:0] taps4x = sub_wire9[804:644];

	altshift_taps	ALTSHIFT_TAPS_component (
				.aclr (aclr),
				.clock (clock),
				.shiftin (shiftin),
				.shiftout (sub_wire0),
				.taps (sub_wire1)
				// synopsys translate_off
				,
				.clken (),
				.sclr ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Cyclone IV GX",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=M9K",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 5,
		ALTSHIFT_TAPS_component.tap_distance = 10,
		ALTSHIFT_TAPS_component.width = 161;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "1"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "5"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "10"
// Retrieval info: PRIVATE: WIDTH NUMERIC "161"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M9K"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "5"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "10"
// Retrieval info: CONSTANT: WIDTH NUMERIC "161"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT VCC "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 161 0 INPUT NODEFVAL "shiftin[160..0]"
// Retrieval info: USED_PORT: shiftout 0 0 161 0 OUTPUT NODEFVAL "shiftout[160..0]"
// Retrieval info: USED_PORT: taps0x 0 0 161 0 OUTPUT NODEFVAL "taps0x[160..0]"
// Retrieval info: USED_PORT: taps1x 0 0 161 0 OUTPUT NODEFVAL "taps1x[160..0]"
// Retrieval info: USED_PORT: taps2x 0 0 161 0 OUTPUT NODEFVAL "taps2x[160..0]"
// Retrieval info: USED_PORT: taps3x 0 0 161 0 OUTPUT NODEFVAL "taps3x[160..0]"
// Retrieval info: USED_PORT: taps4x 0 0 161 0 OUTPUT NODEFVAL "taps4x[160..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 161 0 shiftin 0 0 161 0
// Retrieval info: CONNECT: shiftout 0 0 161 0 @shiftout 0 0 161 0
// Retrieval info: CONNECT: taps0x 0 0 161 0 @taps 0 0 161 0
// Retrieval info: CONNECT: taps1x 0 0 161 0 @taps 0 0 161 161
// Retrieval info: CONNECT: taps2x 0 0 161 0 @taps 0 0 161 322
// Retrieval info: CONNECT: taps3x 0 0 161 0 @taps 0 0 161 483
// Retrieval info: CONNECT: taps4x 0 0 161 0 @taps 0 0 161 644
// Retrieval info: GEN_FILE: TYPE_NORMAL shift.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL shift.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shift.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shift.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shift_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL shift_bb.v TRUE
